//////////////////////////
//
//
//文件名：decode.v
//模块名：DECODE
//创建日期：2022-7-22
//最后修改日期: 2022-7-22
//解码
//
//
//////////////////////////


module DECODE(
    input clk,
    input [31:0] inst,
    output decode_out//TODO: 信号定义
);


endmodule