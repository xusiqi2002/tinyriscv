//////////////////////////
//
//
//文件名：regfile.v
//模块名：RF
//寄存器堆
//此处仅考虑32个通用寄存器
//
//
//创建日期：2022-7-22
//最后修改日期: 2022-7-22
//
//
//////////////////////////
module RF(

);


endmodule